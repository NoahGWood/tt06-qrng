VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO H_WG
  CLASS BLOCK ;
  FOREIGN H_WG ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.010 BY 0.010 ;
END H_WG
END LIBRARY

