magic
tech sky130A-GDS
timestamp 1709357108
<< POLY >>
rect -1 -1 15992 9996
<< end >>
